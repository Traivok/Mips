module TestModule(input logic [31:0] a, 
				  output logic [31:0] b,
				  input logic clk, res, lod);
	Registrador(clk, res, lod, a, b);
endmodule : TestModule