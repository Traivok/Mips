module MIPS(input logic in, output logic out);
	TestModule(in, out);
endmodule : MIPS